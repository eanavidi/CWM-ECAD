//////////////////////////////////////////////////////////////////////////////////
// Exercise #2 - Doorbell Chime
// Student Name:
// Date: 
//
//  Description: In this exercise, you need to design a multiplexer that chooses between two sounds, where the  
//  output is delayed by 5 ticks (not clocks!) and acts according to the following truth table:
//
//  sel | out
// -----------------
//   0  | a
//   1  | b
//
//  inputs:
//           a, b, sel
//
//  outputs:
//           out
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

module MUX(
    input [24:0] a,
    input [24:0] b,
    input sel,
    output reg [24:0] out
    );
  

always @ (*) begin
    #5;
   
       if (sel)
           out = b;

       else
           out = a;
    
end 

endmodule
  
